library verilog;
use verilog.vl_types.all;
entity fourBitComparator_vlg_vec_tst is
end fourBitComparator_vlg_vec_tst;
